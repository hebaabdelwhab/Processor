----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Decoder is
end Decoder;

architecture Behavioral of Decoder is

begin


end Behavioral;

